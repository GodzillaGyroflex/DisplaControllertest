`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:24:05 03/15/2017 
// Design Name: 
// Module Name:    Counter 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

module nBitCounter(count, enable, clk, rst_n);
  parameter n = 15;
 
  output reg [n:0] count;
  input clk;
  input rst_n;
  input enable;
 
  // Set the initial value
  initial
    count = 0;
 
  // Increment count on clock
  always @(posedge clk or negedge rst_n)  
    if (!rst_n)
      count = 0;		
    else if(enable)
      count = count + 1;
	
endmodule

		


